package Regs;

import GetPut::*;
import ClientServer::*;
import RegCommon::*;







endpackage