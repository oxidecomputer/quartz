package Sequencer;

endpackage
